program tb_vm(output bit valid_s,
			  output bit [2:0] items_s,
			  output bit [3:0] count_s,
			  output bit [7:0] cost_s,
			  output bit enter_key,
			  output bit clk,rst,
			  output bit [1:0]coins,
			  output bit [5:0]button,
			  input logic [2:0]product,
              input logic [1:0]status,
              input logic [15:0]balance,
              input logic [7:0]info, 
			  output bit soft_rst
			  );
			  
/*//SUPPLIER INPUTS TO DESIGN
bit valid_s;
bit [2:0] item_s;
bit [3:0] count_s;
bit [7:0] cost_s;
bit enter_key;

//USER INPUTS TO DESIGN
bit [1:0]coins;
bit [5:0]button;

//ESSENTIAL INPUTS
bit clk, rst;*/

//======================= Clock Generator =================================================

initial begin: clockGenerator
	clk = 0;							//Initializing the clk to 0.
	forever #5 clk = ~clk;				//Toggling the clk after every 5 unit time.
end: clockGenerator

//======================== SUPPLIER Task to perform Restocking ============================
task supplier;
		int i;
		valid_s = 1'b1;
		rst = 1'b0;
		for(i=0;i<6;i++)
			begin
				items_s = i;
				cost_s = i*5+5;
				count_s = 15;
			$display("ITEM = %d\t COST = %b\t COUNT =%d",items_s,cost_s,count_s);
				#10;
			end
		valid_s = 1'b0;
endtask: supplier


task buttoncoinzero;
		button = 6'b000000;
		coins = 2'b00;
endtask:buttoncoinzero


task consumer(
			input logic [5:0]i,
			input logic [1:0]j,
			input logic k);
		begin
		//@(posedge clk);
			button = i;
			coins = j;
			enter_key = k;
			
			repeat(2) @(posedge clk)buttoncoinzero;
			#10;
		
				
		end
endtask

//Task for when user putting coins continously.  
task coins_continue(
					input logic [5:0]i,
					input logic [1:0]j,
					input logic k
					);
		begin
			button = i;
			coins = j;
			enter_key = k;
			#10;
		end
endtask:coins_continue

initial
	begin
		$monitor("STATUS=%d\t BUTTON=%b\t COINS=%b\t PRODUCT=%d\t BALANCE =%d\t INFORMATION = %d\t",status,button,coins,product,balance,info);
		
			@(posedge clk)supplier;
//========================= Test Case 1: CONSUMER : BUTTON 1 is SELECTED : COIN 5 cent is inserted ===========================	
			#10 repeat(3) @(posedge clk) consumer(6'b000100,2'b01,1'b1);
			
//========================= Test Case 2: CONSUMER : BUTTON 2 is SELECTED : COIN 5 cent is inserted for 10 cent product value ================
			#10 repeat(2) @(posedge clk) consumer(6'b000010,2'b01,1'b1);
			
//========================= Test Case 3: CONSUMER : BUTTON 2 is SELECTED : COIN 10 cent is inserted continously for 10 cent product value ================			
			#10 repeat(3) @(posedge clk) coins_continue(6'b010000,2'b11,1'b1);
			
//========================= Test Case 4: CONSUMER : BUTTON 1 and 3 is SELECTED : COIN 5 cent is inserted =========================== 	
			#20  @(posedge clk) consumer(6'b000101,2'b01,1'b1);
				
			#200 $stop;
	end
endprogram		
